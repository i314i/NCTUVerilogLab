`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:58:52 10/02/2015 
// Design Name: 
// Module Name:    RING_COUNTER 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RING_COUNTER(
    input clk,
    input rst,
    output reg t0,
	 output reg t1,
	 output reg t2,
	 output reg t3
    );


endmodule
